`ifndef NICE_PATTERNS_TYPEDEFS_SVH
`define NICE_PATTERNS_TYPEDEFS_SVH

typedef interface class iterable;
typedef interface class iterator;
typedef interface class composite;

typedef class enum_iterator;
typedef class composition_iterator;

typedef class composition_leaf;
typedef class composition_node;

typedef class singleton_proxy;


`endif // NICE_PATTERNS_TYPEDEFS_SVH
