//-----------------------------------------------------------------------------
// Project       : Callisto
//-----------------------------------------------------------------------------
// File          : nice_io_types.svh
// Author        : skimhi
// Created       : Mon Sep 2024, 11:22:25
// Last modified : Mon Sep 2024, 11:22:25
//
//-----------------------------------------------------------------------------
// Copyright (c) Speedata.
//------------------------------------------------------------------------------
// Modification history:
// Mon Sep 2024, 11:22:25
//-----------------------------------------------------------------------------

`ifndef NICE_IO_TYPES_SVH
`define NICE_IO_TYPES_SVH

typedef interface class stream;

typedef class file;
typedef class file_reader;
typedef class cmdline_arg;

`endif // NICE_IO_TYPES_SVH
