//-----------------------------------------------------------------------------
// Project       : Callisto
//-----------------------------------------------------------------------------
// File          : nice_patterns_typedefs.svh
// Author        : skimhi
// Created       : Sat Sep 2024, 21:59:41
// Last modified : Sat Sep 2024, 21:59:41
//
//-----------------------------------------------------------------------------
// Copyright (c) Speedata.
//------------------------------------------------------------------------------
// Modification history:
// Sat Sep 2024, 21:59:41
//-----------------------------------------------------------------------------

`ifndef NICE_PATTERNS_TYPEDEFS_SVH
`define NICE_PATTERNS_TYPEDEFS_SVH

typedef interface class iterable;
typedef interface class iterator;
typedef interface class composite;

typedef class enum_iterator;
typedef class composition_iterator;

typedef class composition_leaf;
typedef class composition_node;

typedef class singleton_proxy;


`endif // NICE_PATTERNS_TYPEDEFS_SVH
