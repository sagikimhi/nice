`ifndef NICE_IO_TYPES_SVH
`define NICE_IO_TYPES_SVH

typedef class file;
typedef class file_reader;
typedef class cmdline_arg;
typedef interface class stream;

`endif // NICE_IO_TYPES_SVH
